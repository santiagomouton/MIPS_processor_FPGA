`timescale 1ns / 1ps

module decode_top
	#(
		parameter NB_DATA   = 32,		
		parameter NB_OPCODE = 6,
		parameter NB_REG    = 5				
	)
	(
		input wire clock_i,
		input wire reset_i,
		input wire [7-1:0] pc_decode,
		//input wire enable_i,
		input wire reg_write_i,
		input wire select_debug_or_wireA,	
		input wire [NB_REG-1:0] addr_reg_debug,	
		
		input wire [NB_DATA-1:0] instruction_i,		
		input wire [NB_REG-1:0] write_register_i,
		input wire [NB_DATA-1:0] data_rw_i,

		input wire decode_forward_A, 
        input wire decode_forward_B,
		input wire [NB_DATA-1:0] alu_result,

		input wire stall,

		// output wire [NB_REG-1:0] shamt_o,
		output wire [NB_REG-1:0] wireA_o, wireB_o, wireRW_o,

		output wire [5:0]mem_signals, 
		output wire [2:0]wb_signals,
        output wire [1:0]regDest_signal,
        output wire tipeI_signal,
        output wire shamt_signal,

        output wire [NB_OPCODE-1:0] opcode_o,
        output wire [5:0] funct_o,
        output wire [NB_DATA-1:0] wire_inmediate_sign_o,
        output wire [NB_DATA-1:0] data_ra_o,
        output wire [NB_DATA-1:0] data_rb_o,

		output wire pc_branch_or_jump,
		output wire [7-1:0] address_jump,
		output wire [7-1:0] address_branch,
		output wire [7-1:0] address_register,
		output wire [1:0] pc_src,
		output wire halt_signal,
		output wire [31:0] wire_inmediate_paraver
	);

	wire [NB_REG-1:0] addr_A_out;

	// Conexion distribuidor, banco de registros y control unit
	wire [5:0]operation;
	wire [5:0]funct;
	wire is_equal;

	//distributor
	wire [NB_REG-1:0] wire_A;
	wire [NB_REG-1:0] wire_B;
	wire [26-1:0] wire_direction;
	wire [16-1:0] wire_inmediate;

	// control_unit
	wire [5:0]mem_signals_ctr; 
	wire [2:0]wb_signals_ctr;
	wire [1:0]regDest_signal_ctr;
	wire tipeI_signal_ctr;
	wire beq, bne, jump;
	wire shamt_signal_ctr;
	wire [NB_OPCODE-1:0] opcode_ctr;

	wire [NB_DATA-1:0] data_ra, data_rb, data_ra_branch, data_rb_branch;

	wire [NB_DATA-1:0] wire_inmediate_sign;

	assign data_ra_o = data_ra;
	assign data_rb_o = data_rb;

    assign wireA_o = wire_A;
    assign wireB_o = wire_B;
    // assign funct_o = funct;
	assign wire_inmediate_sign_o = wire_inmediate_sign;

	assign pc_branch_or_jump = ((is_equal && beq) | (!is_equal && bne) | jump);
	assign address_jump 	 = pc_decode + wire_direction[7-1:0]; //acotado porque tomamos solo 32 direcciones de instrucciones en este tp
	assign address_register  = data_ra[7-1:0];

    assign mem_signals 	  = (stall) ? {6'b0} : mem_signals_ctr;
	assign wb_signals     = (stall) ? {3'b0} : wb_signals_ctr;
	assign regDest_signal = (stall) ? {2'b0} : regDest_signal_ctr;
	assign opcode_o 	  = (stall) ? {6'b0} : opcode_ctr;
	assign funct_o 		  = (stall) ? {6'b0} : funct;
	assign tipeI_signal   = (stall) ? (1'b1) : tipeI_signal_ctr;
	assign shamt_signal   = (stall) ? (1'b0) : shamt_signal_ctr;


	branch branch
	(
		.pc(pc_decode),
		.inmediate(wire_inmediate_sign),
		.data_ra_branch(data_ra_branch),
		.data_rb_branch(data_rb_branch),

		.is_equal(is_equal),
		.branch_address_o(address_branch)
	);

 	multiplexor_2_in #(.NB_DATA(NB_REG)) addr_debug_or_wireA
	(
		.op1_i(wire_A),
		.op2_i(addr_reg_debug),
		.sel_i(select_debug_or_wireA),
		.data_o(addr_A_out)
	);

	bank_registers bank_registers
	(
		.clock_i(clock_i),
		.reset_i(reset_i),
		.rw_i(reg_write_i), 
		.addr_ra_i(addr_A_out),
		.addr_rb_i(wire_B),
		.addr_rw_i(write_register_i),
		.data_rw_i(data_rw_i),
		.data_ra_o(data_ra),
		.data_rb_o(data_rb)		
	);
	
	distributor distributor
	(
		.instruction(instruction_i),
		// .regDst(1'b0),
		.operation(operation),
		.funct(funct),
		.inmediate(wire_inmediate),
		.wire_A(wire_A),
		.wire_B(wire_B),
		.direction(wire_direction),
		.wire_dest(wireRW_o)
	);
	assign wire_inmediate_paraver = {16'b0, wire_inmediate};

	control_unit control_unit
	(
        .opcode(operation),
        // .funct(funct),
        .wb_signals(wb_signals_ctr),
		.tipeI(tipeI_signal_ctr),
		
		.shamt(shamt_signal_ctr),
        .beq(beq),
		.bne(bne),
		.jump(jump),
		.pc_src(pc_src),

        .regDest_signal(regDest_signal_ctr),
		.opcode_o(opcode_ctr),
        .mem_signals(mem_signals_ctr),
		.halt_signal(halt_signal)
	);

	sign_extension sign_extension
	(
		.unextend_i(wire_inmediate),
        .extended_o(wire_inmediate_sign) 
	);	

 //OJO CON ESTO, SELECCION QUIZAS INCORRECTA
 	multiplexor_2_in#(.NB_DATA(NB_DATA)) forward_or_reg_A
	(
		.op1_i(data_ra),
		.op2_i(alu_result), //1
		.sel_i(decode_forward_A),
		.data_o(data_ra_branch)
	);
    multiplexor_2_in#(.NB_DATA(NB_DATA)) forward_or_reg_B
	(
		.op1_i(data_rb),
		.op2_i(alu_result),
		.sel_i(decode_forward_B),
		.data_o(data_rb_branch)
	);

endmodule

